parameter Nrows   = 798 ;
parameter Ncol    = 532 ;
